library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.Common.all;

entity IrisDataManager is
	port (
		CLK					:	in		std_logic;
		SelectDataType		:	in		std_logic;
		SelectDataIndex		:	in		unsigned(6 downto 0);
		SelectDataOut		:	out	DataAttributes
	);
end entity IrisDataManager;

architecture arch of IrisDataManager is
	constant TrainingCount	:	integer	:= 120;
	constant TestCount		:	integer	:= 30;
	
	type TrainingDataArray is array(0 to TrainingCount - 1) of DataAttributes;
	type TestDataArray is array(0 to TestCount - 1) of DataAttributes;
	
	-- data set from https://archive.ics.uci.edu/ml/datasets/iris
	-- contains 40 of each class, totaling 120 = 80% of total data set
	-- 1. sepal length in cm
	-- 2. sepal width in cm
	-- 3. petal length in cm
	-- 4. petal width in cm
	-- 5. class:
	--   0.0 -> Iris Setosa
	--   1.0 -> Iris Versicolour
	--   2.0 -> Iris Virginica
	constant TrainingData : TrainingDataArray := (
		(51,35,14,2,0),
		(49,30,14,2,0),
		(47,32,13,2,0),
		(46,31,15,2,0),
		(50,36,14,2,0),
		(54,39,17,4,0),
		(46,34,14,3,0),
		(50,34,15,2,0),
		(44,29,14,2,0),
		(49,31,15,1,0),
		(54,37,15,2,0),
		(48,34,16,2,0),
		(48,30,14,1,0),
		(43,30,11,1,0),
		(58,40,12,2,0),
		(57,44,15,4,0),
		(54,39,13,4,0),
		(51,35,14,3,0),
		(57,38,17,3,0),
		(51,38,15,3,0),
		(54,34,17,2,0),
		(51,37,15,4,0),
		(46,36,10,2,0),
		(51,33,17,5,0),
		(48,34,19,2,0),
		(50,30,16,2,0),
		(50,34,16,4,0),
		(52,35,15,2,0),
		(52,34,14,2,0),
		(47,32,16,2,0),
		(48,31,16,2,0),
		(54,34,15,4,0),
		(52,41,15,1,0),
		(55,42,14,2,0),
		(49,31,15,2,0),
		(50,32,12,2,0),
		(55,35,13,2,0),
		(49,36,14,1,0),
		(44,30,13,2,0),
		(51,34,15,2,0),
		(70,32,47,14,1),
		(64,32,45,15,1),
		(69,31,49,15,1),
		(55,23,40,13,1),
		(65,28,46,15,1),
		(57,28,45,13,1),
		(63,33,47,16,1),
		(49,24,33,10,1),
		(66,29,46,13,1),
		(52,27,39,14,1),
		(50,20,35,10,1),
		(59,30,42,15,1),
		(60,22,40,10,1),
		(61,29,47,14,1),
		(56,29,36,13,1),
		(67,31,44,14,1),
		(56,30,45,15,1),
		(58,27,41,10,1),
		(62,22,45,15,1),
		(56,25,39,11,1),
		(59,32,48,18,1),
		(61,28,40,13,1),
		(63,25,49,15,1),
		(61,28,47,12,1),
		(64,29,43,13,1),
		(66,30,44,14,1),
		(68,28,48,14,1),
		(67,30,50,17,1),
		(60,29,45,15,1),
		(57,26,35,10,1),
		(55,24,38,11,1),
		(55,24,37,10,1),
		(58,27,39,12,1),
		(60,27,51,16,1),
		(54,30,45,15,1),
		(60,34,45,16,1),
		(67,31,47,15,1),
		(63,23,44,13,1),
		(56,30,41,13,1),
		(55,25,40,13,1),
		(63,33,60,25,2),
		(58,27,51,19,2),
		(71,30,59,21,2),
		(63,29,56,18,2),
		(65,30,58,22,2),
		(76,30,66,21,2),
		(49,25,45,17,2),
		(73,29,63,18,2),
		(67,25,58,18,2),
		(72,36,61,25,2),
		(65,32,51,20,2),
		(64,27,53,19,2),
		(68,30,55,21,2),
		(57,25,50,20,2),
		(58,28,51,24,2),
		(64,32,53,23,2),
		(65,30,55,18,2),
		(77,38,67,22,2),
		(77,26,69,23,2),
		(60,22,50,15,2),
		(69,32,57,23,2),
		(56,28,49,20,2),
		(77,28,67,20,2),
		(63,27,49,18,2),
		(67,33,57,21,2),
		(72,32,60,18,2),
		(62,28,48,18,2),
		(61,30,49,18,2),
		(64,28,56,21,2),
		(72,30,58,16,2),
		(74,28,61,19,2),
		(79,38,64,20,2),
		(64,28,56,22,2),
		(63,28,51,15,2),
		(61,26,56,14,2),
		(77,30,61,23,2),
		(63,34,56,24,2),
		(64,31,55,18,2),
		(60,30,48,18,2),
		(69,31,54,21,2)
	);
	
	-- contains 10 of each class, totaling 30 = 20% of total data set
	constant TestData : TestDataArray := (
		(50,35,13,3,0),
		(45,23,13,3,0),
		(44,32,13,2,0),
		(50,35,16,6,0),
		(51,38,19,4,0),
		(48,30,14,3,0),
		(51,38,16,2,0),
		(46,32,14,2,0),
		(53,37,15,2,0),
		(50,33,14,2,0),
		(55,26,44,12,1),
		(61,30,46,14,1),
		(58,26,40,12,1),
		(50,23,33,10,1),
		(56,27,42,13,1),
		(57,30,42,12,1),
		(57,29,42,13,1),
		(62,29,43,13,1),
		(51,25,30,11,1),
		(57,28,41,13,1),
		(67,31,56,24,2),
		(69,31,51,23,2),
		(58,27,51,19,2),
		(68,32,59,23,2),
		(67,33,57,25,2),
		(67,30,52,23,2),
		(63,25,50,19,2),
		(65,30,52,20,2),
		(62,34,54,23,2),
		(59,30,51,18,2)	
	);

	constant NullData : DataAttributes := (0, 0, 0, 0, 0);
begin
	process(CLK)
	begin
		if (CLK'event and CLK = '1') then
			if (SelectDataType = '0') then
				SelectDataOut <= TrainingData(to_integer(SelectDataIndex));
			elsif (SelectDataType = '1') then
				SelectDataOut <= TestData(to_integer(SelectDataIndex));
			else
				SelectDataOut <= NullData;
			end if;
		end if;
	end process;
end architecture arch;